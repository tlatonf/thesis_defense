`define B_WIDTH     1600
`define W_WIDTH     64
`define L_WIDTH     6

`define C_WIDTH     1024
`define R_WIDTH     576

`define NR          24  // Number of rounds

`define ENABLE      1'b1
`define DISABLE     1'b0

`define TYPE_SHA3_512   2'b00
`define TYPE_SHA3_256   2'b01
`define TYPE_SHAKE_128  2'b10
`define TYPE_SHAKE_256  2'b11