function logic [0:63] rot;
  // rotate left
  input logic [0:63] in;
  input logic [0:5] n;
  begin
    case (n)
      6'd0:  rot = in;
      6'd1:  rot = {in[ 1:63], in[0   ]};
      6'd2:  rot = {in[ 2:63], in[0: 1]};
      6'd3:  rot = {in[ 3:63], in[0: 2]};
      6'd4:  rot = {in[ 4:63], in[0: 3]};
      6'd5:  rot = {in[ 5:63], in[0: 4]};
      6'd6:  rot = {in[ 6:63], in[0: 5]};
      6'd7:  rot = {in[ 7:63], in[0: 6]};
      6'd8:  rot = {in[ 8:63], in[0: 7]};
      6'd9:  rot = {in[ 9:63], in[0: 8]};
      6'd10: rot = {in[10:63], in[0: 9]};
      6'd11: rot = {in[11:63], in[0:10]};
      6'd12: rot = {in[12:63], in[0:11]};
      6'd13: rot = {in[13:63], in[0:12]};
      6'd14: rot = {in[14:63], in[0:13]};
      6'd15: rot = {in[15:63], in[0:14]};
      6'd16: rot = {in[16:63], in[0:15]};
      6'd17: rot = {in[17:63], in[0:16]};
      6'd18: rot = {in[18:63], in[0:17]};
      6'd19: rot = {in[19:63], in[0:18]};
      6'd20: rot = {in[20:63], in[0:19]};
      6'd21: rot = {in[21:63], in[0:20]};
      6'd22: rot = {in[22:63], in[0:21]};
      6'd23: rot = {in[23:63], in[0:22]};
      6'd24: rot = {in[24:63], in[0:23]};
      6'd25: rot = {in[25:63], in[0:24]};
      6'd26: rot = {in[26:63], in[0:25]};
      6'd27: rot = {in[27:63], in[0:26]};
      6'd28: rot = {in[28:63], in[0:27]};
      6'd29: rot = {in[29:63], in[0:28]};
      6'd30: rot = {in[30:63], in[0:29]};
      6'd31: rot = {in[31:63], in[0:30]};
      6'd32: rot = {in[32:63], in[0:31]};
      6'd33: rot = {in[33:63], in[0:32]};
      6'd34: rot = {in[34:63], in[0:33]};
      6'd35: rot = {in[35:63], in[0:34]};
      6'd36: rot = {in[36:63], in[0:35]};
      6'd37: rot = {in[37:63], in[0:36]};
      6'd38: rot = {in[38:63], in[0:37]};
      6'd39: rot = {in[39:63], in[0:38]};
      6'd40: rot = {in[40:63], in[0:39]};
      6'd41: rot = {in[41:63], in[0:40]};
      6'd42: rot = {in[42:63], in[0:41]};
      6'd43: rot = {in[43:63], in[0:42]};
      6'd44: rot = {in[44:63], in[0:43]};
      6'd45: rot = {in[45:63], in[0:44]};
      6'd46: rot = {in[46:63], in[0:45]};
      6'd47: rot = {in[47:63], in[0:46]};
      6'd48: rot = {in[48:63], in[0:47]};
      6'd49: rot = {in[49:63], in[0:48]};
      6'd50: rot = {in[50:63], in[0:49]};
      6'd51: rot = {in[51:63], in[0:50]};
      6'd52: rot = {in[52:63], in[0:51]};
      6'd53: rot = {in[53:63], in[0:52]};
      6'd54: rot = {in[54:63], in[0:53]};
      6'd55: rot = {in[55:63], in[0:54]};
      6'd56: rot = {in[56:63], in[0:55]};
      6'd57: rot = {in[57:63], in[0:56]};
      6'd58: rot = {in[58:63], in[0:57]};
      6'd59: rot = {in[59:63], in[0:58]};
      6'd60: rot = {in[60:63], in[0:59]};
      6'd61: rot = {in[61:63], in[0:60]};
      6'd62: rot = {in[62:63], in[0:61]};
      6'd63: rot = {in[63   ], in[0:62]};
    endcase      
  end
endfunction

function logic [0:63] get_rc;
  input logic [0:4] ir;
  begin
    case (ir)
      5'd0 : get_rc = 64'h0000000000000001;
      5'd1 : get_rc = 64'h0000000000008082;
      5'd2 : get_rc = 64'h800000000000808A;
      5'd3 : get_rc = 64'h8000000080008000;
      5'd4 : get_rc = 64'h000000000000808B;
      5'd5 : get_rc = 64'h0000000080000001;
      5'd6 : get_rc = 64'h8000000080008081;
      5'd7 : get_rc = 64'h8000000000008009;
      5'd8 : get_rc = 64'h000000000000008A;
      5'd9 : get_rc = 64'h0000000000000088;
      5'd10: get_rc = 64'h0000000080008009;
      5'd11: get_rc = 64'h000000008000000A;
      5'd12: get_rc = 64'h000000008000808B;
      5'd13: get_rc = 64'h800000000000008B;
      5'd14: get_rc = 64'h8000000000008089;
      5'd15: get_rc = 64'h8000000000008003;
      5'd16: get_rc = 64'h8000000000008002;
      5'd17: get_rc = 64'h8000000000000080;
      5'd18: get_rc = 64'h000000000000800A;
      5'd19: get_rc = 64'h800000008000000A;
      5'd20: get_rc = 64'h8000000080008081;
      5'd21: get_rc = 64'h8000000000008080;
      5'd22: get_rc = 64'h0000000080000001;
      5'd23: get_rc = 64'h8000000080008008;
      default: get_rc = 64'h0000000000000000;
    endcase
  end
endfunction